module bug (
    inout wire gpio
);

endmodule
