module top(
	inout x,
	input a
);

assign x = a;

endmodule